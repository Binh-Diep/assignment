module decoder4to16(
    //inputs
    input logic [3:0] x_i,
    //outputs
    output logic [15:0] y_i
);
    //code
    always_comb begin
        case (x_i[3:0])
            4'b0000: y_i = 16'b1000000000000000;
            4'b0001: y_i = 16'b0100000000000000; 
            4'b0010: y_i = 16'b0010000000000000; 
            4'b0011: y_i = 16'b0001000000000000; 
            4'b0100: y_i = 16'b0000100000000000; 
            4'b0101: y_i = 16'b0000010000000000; 
            4'b0110: y_i = 16'b0000001000000000; 
            4'b0111: y_i = 16'b0000000100000000;
            4'b1000: y_i = 16'b0000000010000000;
            4'b1001: y_i = 16'b0000000001000000;
            4'b1010: y_i = 16'b0000000000100000;
            4'b1011: y_i = 16'b0000000000010000;
            4'b1100: y_i = 16'b0000000000001000;
            4'b1101: y_i = 16'b0000000000000100;
            4'b1110: y_i = 16'b0000000000000010;
            4'b1111: y_i = 16'b0000000000000001;
            default: y_i = 16'h0;
        endcase
    end
endmodule : decoder4to16
