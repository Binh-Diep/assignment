module encoder16to4(
    //inputs
    input logic [15:0] x_i,
    //outputs
    output logic [3:0] y_i
);
    //code
    always_comb begin
        casez (x_i[15:0])
            16'b1???????????????: y_i = 4'b0000;
            16'b01??????????????: y_i = 4'b0001;
            16'b001?????????????: y_i = 4'b0010;
            16'b0001????????????: y_i = 4'b0011;
            16'b00001???????????: y_i = 4'b0100;
            16'b000001??????????: y_i = 4'b0101;
            16'b0000001?????????: y_i = 4'b0110;
            16'b00000001????????: y_i = 4'b0111;
            16'b000000001???????: y_i = 4'b1000;
            16'b0000000001??????: y_i = 4'b1001;
            16'b00000000001?????: y_i = 4'b1010;
            16'b000000000001????: y_i = 4'b1011;
            16'b0000000000001???: y_i = 4'b1100;
            16'b00000000000001??: y_i = 4'b1101;
            16'b000000000000001?: y_i = 4'b1110;
            16'b0000000000000001: y_i = 4'b1111;
            default: y_i = 4'b0000;
        endcase
    end
endmodule : encoder16to4
